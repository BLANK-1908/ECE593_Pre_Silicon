typedef enum {and_op,exor_op,add_op,mul_op,store_op,load_op} opcodes;
