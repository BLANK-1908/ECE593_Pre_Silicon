
`include "N:/Desktop/Cache/tb.sv" //add your own file directory
`include "N:/Desktop/Cache/top.sv"
