
package filepackage;

`include "packet.sv"

endpackage