`include "tb.sv"
`include "top.sv"
